LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECOFIN IS
	PORT(NUM: IN INTEGER RANGE 1 TO 5; 
			  S1, S2, S3, S4, S5: OUT STD_LOGIC); -- PARA LOS 8 SEG DEL DISPLAY
END ENTITY;

ARCHITECTURE BEAS OF DECOFIN IS
BEGIN
	PROCESS(NUM)
	BEGIN
			IF NUM=1 THEN
				S1<='0';
			ELSIF NUM=2 THEN
				S2<='0';
			ELSIF NUM=3 THEN
				S3<='0';
			ELSIF NUM=4 THEN
				S4<='0';
			ELSE 
				S5<='0';
			END IF;
	END PROCESS;
END BEAS;
