LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY decc IS
	PORT(	R: IN INTEGER RANGE 0 TO 999;
			U, D, C: OUT INTEGER RANGE 0 TO 10);
			
END ENTITY;

ARCHITECTURE BEAS OF decc IS
BEGIN
	
			U<=R MOD 10;
			D<=(R/10) MOD 10;
			C<= (R/100) MOD 10;

END BEAS;