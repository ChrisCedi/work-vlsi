LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM2 IS
	PORT(CLK: IN STD_LOGIC;
			R, ENT: IN INTEGER RANGE 0 TO 999;
			L: OUT INTEGER RANGE 1 TO 3;
			WL: OUT INTEGER RANGE 4 TO 5;
			REINICIA: OUT STD_LOGIC;
			TIEMPO: OUT INTEGER RANGE 1 TO 5);
END ENTITY;

ARCHITECTURE BEAS OF FSM2 IS
TYPE EDOS IS (INI, E1, WIN, LOSE);
SIGNAL LEVEL : INTEGER RANGE 1 TO 3 := 1;
SIGNAL PRES: EDOS := INI;
BEGIN

	PROCESS(R, ENT, CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			CASE PRES IS
				WHEN INI =>
					L <= LEVEL;
					PRES <= E1;
				WHEN E1 => 
					IF LEVEL = 3 THEN
						PRES <= WIN;
					ELSE
						IF R = ENT THEN
							LEVEL <= LEVEL + 1;
							REINICIA <= '1';
							PRES <= INI;
						ELSE
							PRES <= LOSE;
						END IF;
					END IF;
					
				WHEN WIN =>
					WL <= 4;
					
				WHEN LOSE =>
					WL <= 5;
				
			END CASE;
		END IF;
	END PROCESS;

END BEAS;