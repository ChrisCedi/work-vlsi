LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DECASC IS
    PORT (
        ASCCI : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        NUM: OUT INTEGER RANGE 0 TO 9);
		  
END ENTITY;

ARCHITECTURE BEAS OF DECASC IS
BEGIN
    PROCESS(ASCCI)
	 BEGIN
        CASE ASCCI IS
            WHEN "00110000" => NUM <= 0; 
            WHEN "00110001" => NUM <= 1; 
            WHEN "00110010" => NUM <= 2; 
            WHEN "00110011" => NUM <= 3; 
            WHEN "00110100" => NUM <= 4; 
            WHEN "00110101" => NUM <= 5; 
            WHEN "00110110" => NUM <= 6; 
            WHEN "00110111" => NUM <= 7; 
            WHEN "00111000" => NUM <= 8; 
            WHEN "00111001" => NUM <= 9; 
            WHEN OTHERS => NUM <= 0; 
        END CASE;
    END PROCESS;
END BEAS;

