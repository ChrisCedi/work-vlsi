LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY UNIR IS
	PORT(	DIG: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			ENT: OUT STD_LOGIC_VECTOR(9 DOWNTO 0));
END ENTITY;

ARCHITECTURE BEAS OF UNIR IS
BEGIN
END BEAS;