LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SEPAENT IS
	PORT(	R: IN INTEGER RANGE 0 TO 999;
			U2, D2, C2: OUT INTEGER RANGE 0 TO 10);
END ENTITY;

ARCHITECTURE BEAS OF SEPAENT IS
SIGNAL TIEMPO: INTEGER RANGE 0 TO 8 :=0;
BEGIN
	
			U2<=R MOD 10;
			D2<=(R/10) MOD 10;
			C2<= (R/100) MOD 10;

END BEAS;