LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CUAL IS
	PORT(U1, D1, C1: IN INTEGER RANGE 0 TO 10;
			AC: IN STD_LOGIC;
			U2, D2, C2: IN INTEGER RANGE 0 TO 10;
			U, D, C: OUT INTEGER RANGE 0 TO 10);
END ENTITY;

ARCHITECTURE BEAS OF CUAL IS
BEGIN
	PROCESS(AC)
	BEGIN 
		IF AC='1' THEN
			U <= U2;
			D <= D2;
			C <= C2;
		ELSE 
			U <= U1;
			D <= D1;
			C <= C1;
		END IF;
	END PROCESS;
END BEAS;