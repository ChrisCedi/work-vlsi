LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY rx_uart IS
PORT(CLK: IN STD_LOGIC;
      RX: IN STD_LOGIC;
	 DATA: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	 RX_FLAG: BUFFER STD_LOGIC;
	 BUSY: OUT STD_LOGIC);
END rx_uart;

ARCHITECTURE BEAS OF rx_uart IS
SIGNAL INDEX: INTEGER RANGE 0 TO 9 := 0;
SIGNAL PRESCL: INTEGER RANGE 0 TO 434 := 0; -- PARA BAUDAJE PRESCL = 50 MHz/115200
SIGNAL DATA_AUX: STD_LOGIC_VECTOR(9 DOWNTO 0);

BEGIN

	PROCESS(CLK)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			IF (RX_FLAG = '0' AND RX = '0') THEN
				INDEX <= 0; -- INICIAR EN POSICIÓN CERO
				PRESCL <= 0;
				BUSY <= '1'; -- PUERTO SERIE OCUPADO
				RX_FLAG <= '1'; -- ESTA RECIBIENDO
			END IF;
		
			IF RX_FLAG = '1' THEN
				DATA_AUX(INDEX) <= RX;
				IF PRESCL < 434 THEN
					PRESCL <= PRESCL + 1;
				ELSE
					PRESCL <= 0;
				END IF;	
			END IF;
			
			IF PRESCL = 217 THEN
				IF INDEX < 9 THEN
					INDEX <= INDEX + 1;
				ELSE
					IF (DATA_AUX(0) = '0' AND DATA_AUX(9) = '1') THEN -- START = 0 & STOP = 1
						DATA <= DATA_AUX(8 DOWNTO 1);
					ELSE
						DATA <= (OTHERS => '0');
					END IF;
					RX_FLAG <= '0';
					BUSY <= '0';
				END IF;
			END IF;
		END IF;
		
	END PROCESS;
END BEAS;