LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RANDOM IS
	PORT(CLK, STOP: IN STD_LOGIC;
		 AL: OUT INTEGER RANGE 100000000 TO 999999999);
END ENTITY;

ARCHITECTURE BEAS OF RANDOM IS
SIGNAL CUENTA: INTEGER RANGE 100000000 TO 999999999;
BEGIN

	PROCESS(CLK)
	BEGIN
		IF FALLING_EDGE (CLK) THEN
			IF STOP='0' THEN
				AL <= CUENTA;
			ELSE
				IF CUENTA = 999999999 THEN
					CUENTA <= 100000000;
				ELSE
					CUENTA <= CUENTA + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;

END BEAS;